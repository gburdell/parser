`define N 4
