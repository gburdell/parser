`include "./b.vh"
`include "c.vh"

module `MOD ;
	parameter N = `N;
endmodule
