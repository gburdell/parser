`define N 10
