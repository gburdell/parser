`define MOD a
