module foo; i
/* block comment
with //line comment
*/
	"string literal"
input foo; //line comment /*block comment*/
endmodule

	"string which \
	spans multiple lines \"\
	"

	/*block comment with "string"
	*/

