`define M1 4
