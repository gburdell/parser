`include "m1.vh"

module m1; endmodule
